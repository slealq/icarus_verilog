module up_counter_tb {

// initial begin
 input  out;
 output enable;
 output clk;


}
endmodule
